////////

module simple_in_n_out (
    // Inputs
    in_1,
    in_2,
    in_3,
    // Outputs
    out_1,
    out_2
    );

    // Port definition

    input in_1;
    input in_2;
    input in_3;

    output out_1;
    output out_2;

    // Design implementation
    assign out_1 = in_1 & in_2 & in_3;
    assign out_2 = in_1 | in_2 | in_3;
    
endmodule

module intermediate_sig (
    // Inputs
    in_1,
    in_2,
    in_3,
    // Outputs
    out_1,
    out_2
    );

    // Port definitions
    input in_1;
    input in_2;
    input in_3;

    output out_1;
    output out_2;

    // Defino una señal intermedia
    wire intermediate_sig;

    // Design implementation

    assign intermediate_sig = in_1 & in_2;

    assign out_1 = intermediate_sig & in_3;
    assign out_2 = intermediate_sig | in_3;
    
endmodule