module shiftreg (
    output [3:0] o_led,
    input i_valid,
    input i_reset,
    input clock
);
    
endmodule