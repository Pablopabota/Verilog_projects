// 2 input AND gate model
module and2(A, B, Y);
    input A;
    input B;
    output Y;

assign Y = A & B;

endmodule